library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- Libreria para utilizar el operador '+' y la función CONV_INTEGER 
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity REGISTROS is
    GENERIC( NADDR : INTEGER := 4 ;
             NDATA : INTEGER := 16 );

    Port ( 
           
           -- WRITE REGISTER, SELECCIONA UNO DE LOS 16 REGISTROS PARA ESCRIBIR EL DATO ALMACENADO EN WRITE_DATA 
           WRITE_REGISTER  : in  STD_LOGIC_VECTOR (NADDR-1 downto 0); 
           -- READ REGISTER 1, SELECCIONA UNO DE LOS 16 REGISTROS PARA LEER SU CONTENIDO
           READ_REGISTER1 : in STD_LOGIC_VECTOR (NADDR-1 downto 0);
           READ_REGISTER2 : in STD_LOGIC_VECTOR (NADDR-1 downto 0);
           -- REGISTRO CORRIMIENTO, CONTIENE EL NÚMERO DE CORRIMIENTOS QUE SE APLICARÁN A UN DATO (NUM. DE BITS QUE SE VAN A DESPLAZAR, A LA IZQUIERDA O LA DERECHA) 
           SHAMT: in ST_LOGIC_VECTOR (NADDR-1 DOWNTO 0);
           -- SEÑALES DE CONTROL DEL ARCHIVO DE REGISTROS
           WR, CLK: in STD_LOGIC;
           SHE, DIR: in STD_LOGIC;
           -- MEMORIA RAM MULTIPUERTO, EN ESTE CASO TENEMOS 3, LOS CUALES SON LOS SIGUIENTES:
            -- Bus de datos de entrada WRITE DATA, ES ESTE BUS SE ENCUENTRA EL DATO QUE SE ESCRIBIRÁ EN ALGUNO DE LOS 16 REGISTROS
           WRITE_DATA  : in  STD_LOGIC_VECTOR (NDATA-1 downto 0);
           -- Señales de salida del Archivo de registros
           -- READ_DATA1 ES SALIDA Y ENTRADA, PORQUE ESTA SEÑAL SE RETROALIMENTA AL BLOQUE DE BARREL SHIFTER A SU VEZ QUE SALE CON EL VALOR QUE TIENE EL REGISTRO QUE SE LEYO
           READ_DATA1 : inout ST_LOGIC_VECTOR (NDATA-1 DOWNTO 0);
           READ_DATA2 : out ST_LOGIC_VECTOR (NDATA-1 DOWNTO 0);

end REGISTROS;


architecture ARCHIVO of REGISTROS is
    TYPE MEMORIA IS ARRAY ( (2**NADDR)-1 DOWNTO 0) OF STD_LOGIC_VECTOR(WRITE_DATA'RANGE);
    -- R0 ... R15
    SIGNAL REGS : MEMORIA;
    -- SALIDA DEL MULTIPLEXOR QUE TIENE COMO ENTRADAS WRITE_DATA Y LA SALIDA DE BARREL_SHIFTER
    SIGNAL DATA, DATA_SHIFT : STD_LOGIC_VECTOR( WRITE_DATA'RANGE );
    -- DATA_SHIFT ES LA SALIDA DEL BLOQUE LLAMADO 'BARRELL SHIFTER' QUE SE ENCARGA DE REALIZAR CORRIMIENTOS
    begin 
    -- PROGRAMACIÓN DEL BLOQUE BARRELSHIFTER 
    -- LISTA SENSIBLE DEL BARREL SHIFTER IRAN LAS SEÑALES DE ENTRADA DE ESTE BLOQUE, ESTÁS SERÁN READ_DATA1 (ESTA SEÑAL SE RETROALIMENTA AL BLOQUE DE BARREL SHIFTER), TIENE OTRA ENTRADA LLAMADA SHAMT(NÚMERO DE CORRIMIENTOS QUE SE APLICARÁN) 
    -- Y DIR, ESTA ÚLTIMA SEÑAL INDICA LA DIRECCIÓN DEL CORRIMIENTO, YA SEA A LA IZQUIERDA O A LA DERECHA. 
    BARREL: PROCESS( READ_DATA1, SHAMT, DIR)
        begin
            -- INSTRUCCIÓN DE ALTO NIVEL DE VHDL 
            -- OPERACIÓN DE CORRIMIENTO  BITVECTOR <= TIPO-BITVECTOR SRL TIPO-INTEGER
            -- sll desplazamiento lógico a la iquierda, srl desplazamiento lógico a la derecha
            -- señal, operador, número de bits a recorrer, el desplazamiento se rellena con ceros, ya sea a la izquierda o a la derecha
            -- A LA SEÑAL A LA CUAL YO LE APLICO EL CORRIEMIENTO DEBE SER UNA SEÑAL DE TIPO BIT ESPECÍFICAMENTE (YA QUE ASÍ TRABAJAN LAS OPERACIONES SSL Y SRL, CON SEÑALES DE TIPO BIT), 
            -- COMO NOSOTROS TENEMOS STD_LOGIC_VECTOR, NECESITAMOS HACER UNA CONVERSIÓN DE TIPO, PARA QUE PODAMOS UTILIZAR LAS OPERATIONCES DE CORRIMIENTO
            -- PREGUNTAMOS POR EL VALOR DE DIR
            IF( DIR = '0' ) THEN -- DIR 0 = CORRIMIENTO A LA DERECHA
            -- EN LAS OPERACIONES DE CORRIMIENTO EL NÚMERO DE BITS QUE VOY A RECORRER EN ESTE CASO 'SHAMT' EL VALOR DEBE DE SER UN ENTERO, EL NÚMERO DE BITS A RECORRER DEBE DE SER UN NÚMERO ENTERO
            -- 'INTEGER' POR LO QUE HAREMOS UNA CONVERSIÓN DE TIPO EN SHAMT PARA CONVERTIRLO A UN ENTERO
                DATA_SHIFT <= TO_STDLOGICVECTOR( TO_BITVECTOR(READ_DATA1) SRL CONV_INTEGER(SHAMT) ); -- EL RESULTADO DEL CORRIMIENTO LO PONDREMOS EN DATA_SHIFT
            ELSE 
                -- EL RESULTADO DE UNA OPERACIÓN DE CORRIMIENTO ES DE TIPO BITVECTOR, PERO LO ESTAMOS ASIGNANDO A LA SEÑAL DATA_SHIFT, PERO ESTA ES DE TIPO STD_LOGIC_VECTOR
                -- POR LO QUE HAY QUE HACER OTRA CONVERSIÓN DE TIPO, AHORA CONVERTIREMOS DE BITVECTOR A STD_LOGIC_VECTOR
                DATA_SHIFT <= TO_STDLOGICVECTOR( TO_BITVECTOR(READ_DATA1) SLL CONV_INTEGER(SHAMT) ); -- SI DIR 1 = CORRIMIENTO A LA IZQUIERDA
            END IF;
        end process BARREL;
    -- Programación del multiplexor que tiene como entradas WRITE DATA (CON CERO SE SELECCIONA ESTA) Y DATA_SHIFT (CON UNO DE LA SEÑAL 'SHE' SE LECCIONA ESTA)
    DATA <= WRITE_DATA WHEN ( SHE == '0' ) ELSE DATA_SHIFT;
    -- CUANDO SHE == 0 EN LOS REGISTROS SE ALMACENARÁ EL VALOR QUE TENGA EL BUS WRITE_DATA
    -- CUANDO SHE == 1 EN LOS REGISTROS SE ALMACENARÁ EL VALOR QUE SALGA DEL BLOQUE BARREL_SHIFTER
    
    -- Proceso secuencial
    PMEMDAT : process( CLK )
    -- Proceso de escritura síncrono
    begin       
        IF ( RISING_EDGE(CLK) ) THEN
        -- CUANDO LA SEÑAL WR SEA UNO, SE ESCRIBIRÁ EN ALGUNO DE LOS REGISTROS    
        IF ( WR = '1' ) THEN
                -- EL BUS WRITE REGISTER SELECCIONA EL REGISTRO EN EL QUE YO QUIERO ESCRIBIR
                -- EL VALOR QUE SE VA A ESCRIBIR EN ALGUNO DE LOS REGISTROS ES EL QUE SALE DEL MULTIPLEXOR QUE TIENE COMO ENTRADA WRITE DATA Y LA SALIDA DE BARREL SHIFTER, A ESA SEÑAL DE SALIDA LE LLAMAREMOS 'DATA'
                REGS( CONV_INTEGER(WRITE_REGISTER) ) <= DATA;
            END IF;  
        END IF;
    end process PMEMDAT;
   -- LA LECTURA DE LA MEMORIA ES LA SALIDA DE LOS MULTIPLEXORES, LOS SELECTORES DE CADA 
   -- MULTIPLEXOR SERÁN READ_REGISTER1 y READ_REGISTER2 respectivamente.
    READ_DATA1 <= REGS( CONV_INTEGER(READ_REGISTER1) );
    -- Otro multiplexor de salida.
    READ_DATA2 <= REGS( CONV_INTEGER(READ_REGISTER2) );

end ARCHIVO;